`timescale 1ns / 1ps

//------------------------------------------------------------------------------
// Module: InstROM
// Brief : Instruction memory initialized with sample program words.
//------------------------------------------------------------------------------
module InstROM (
  input  [31:0] Addr,  // Addr-Instruction address
  output [31:0] Inst   // Inst-Instruction
);

  reg [31:0] InstROM[255:0]; // InstROM-Instruction memory

  assign Inst = InstROM[Addr[9:2]];
  integer i;
  initial begin
    for (i = 0; i < 256; i = i + 1) InstROM[i] = 32'h00000000;

    InstROM[0]   = 32'b00110100000000010000000000000101;             // ori $1, $0, 5       # $1 = 5
    InstROM[1]   = 32'b00110100000000100000000000000101;             // ori $2, $0, 5       # $2 = 5
    InstROM[2]   = 32'b00010000001000100000000000000010;             // beq $1, $2, 2       # 相等，跳转到第6行
    InstROM[3]   = 32'b00000000100001010001100000100000;             // add $3, $4, $5      # 不应执行（被冲刷）
    InstROM[4]   = 32'b00000000111010000011000000100010;             // sub $6, $7, $8      # 不应执行（被冲刷）
    InstROM[5]   = 32'b00110100000010010000000000001010;             // ori $9, $0, 10      # 跳转目标，应该执行
    InstROM[6]   = 32'b00110100000010100000000000000001;             // ori $10, $0, 1      # $10 = 1
    InstROM[7]   = 32'b00110100000010110000000000000010;             // ori $11, $0, 2      # $11 = 2
    InstROM[8]   = 32'b00010001010010110000000000000001;             // beq $10, $11, 1     # 不相等，不跳转
    InstROM[9]   = 32'b00000001010010110110000000100000;             // add $12, $10, $11   # 应该执行
    InstROM[10]  = 32'b00110100000011010000000001100100;             // ori $13, $0, 100    # 应该执行
  end
  
endmodule

