`timescale 1ns / 1ps

//------------------------------------------------------------------------------
// Module: InstROM
// Brief : Instruction memory initialized with sample program words.
//------------------------------------------------------------------------------
module InstROM (
  input  [31:0] Addr,  // Addr-Instruction address
  output [31:0] Inst   // Inst-Instruction
);

  reg [31:0] InstROM[255:0]; // InstROM-Instruction memory

  assign Inst = InstROM[Addr[9:2]];
  integer i;
  initial begin
    for (i = 0; i < 256; i = i + 1) InstROM[i] = 32'h00000000;

    // Test program for control hazard handling
    InstROM[0] = 32'b00110100000000010000000000000001;  // ori $1, $0, 1      # $1 = 1
    InstROM[1] = 32'b00110100000000100000000000000010;  // ori $2, $0, 2      # $2 = 2
    InstROM[2] = 32'b00110100000000110000000000000011;  // ori $3, $0, 3      # $3 = 3
    
    // Test BEQ (branch equal) - should not branch
    InstROM[3] = 32'b00010000001000100000000000000010;  // beq $1, $2, 2      # $1 != $2, no branch
    InstROM[4] = 32'b00110100000001000000000000000100;  // ori $4, $0, 4      # $4 = 4 (executed)
    InstROM[5] = 32'b00110100000001010000000000000101;  // ori $5, $0, 5      # $5 = 5 (executed)
    
    // Test BEQ (branch equal) - should branch
    InstROM[6] = 32'b00110100000001100000000000000001;  // ori $6, $0, 1      # $6 = 1
    InstROM[7] = 32'b00010000001001100000000000000010;  // beq $1, $6, 2      # $1 == $6, branch to PC+4+8
    // These two should be flushed:
    InstROM[8] = 32'b00110100000001110000000000000111;  // ori $7, $0, 7      # $7 = 7 (flushed)
    InstROM[9] = 32'b00110100000010000000000000001000;  // ori $8, $0, 8      # $8 = 8 (flushed)
    // Branch target:
    InstROM[10] = 32'b00110100000010010000000000001001; // ori $9, $0, 9      # $9 = 9 (executed)
    
    // Test jump
    InstROM[11] = 32'b00001000000000000000000000001110; // j 14               # Jump to address 14
    // These should be flushed:
    InstROM[12] = 32'b00110100000010100000000000001010; // ori $10, $0, 10    # (flushed)
    InstROM[13] = 32'b00110100000010110000000000001011; // ori $11, $0, 11    # (flushed)
    // Jump target:
    InstROM[14] = 32'b00110100000011000000000000001100; // ori $12, $0, 12    # $12 = 12 (executed)
  end
  
endmodule

