`timescale 1ns / 1ps

//------------------------------------------------------------------------------
// Module: InstROM
// Brief : Instruction memory initialized with sample program words.
//------------------------------------------------------------------------------
module InstROM (
  input  [31:0] Addr,  // Addr-Instruction address
  output [31:0] Inst   // Inst-Instruction
);

  reg [31:0] InstROM[255:0]; // InstROM-Instruction memory

  assign Inst = InstROM[Addr[9:2]];
  integer i;
  initial begin
    for (i = 0; i < 256; i = i + 1) InstROM[i] = 32'h00000000;

    InstROM[0]   = 32'b00000000000000000000000000000000;             // nop
    InstROM[1]   = 32'b10001100000111110000000000000000;             // lw $31, 0($0)
    InstROM[2]   = 32'b00000000000111111111000000100010;             // sub $30, $0, $31
    InstROM[3]   = 32'b00000010000111111110100000100000;             // add $29, $16, $31
    InstROM[4]   = 32'b00000000000111011110000000100010;             // sub $28, $0, $29
    InstROM[5]   = 32'b00000010000111001101100000100000;             // add $27, $16, $28
    InstROM[6]   = 32'b00000011111000011101000000100011;             // subu $26, $31, $1
    InstROM[7]   = 32'b00000000001111111100100000101010;             // slt $25, $1, $31
    InstROM[8]   = 32'b00000000001111111100000000101011;             // sltu $24, $1, $31
    InstROM[9]   = 32'b00100100000101111010101100000000;             // addiu $23, $0, 0xab00
    InstROM[10]  = 32'b00100100000101100000000011001101;             // addiu $22, $0, 0x00cd
    InstROM[11]  = 32'b00110110110101011010101100000000;             // ori $21, $22, 0xab00
    InstROM[12]  = 32'b10101100000101010000000000100000;             // sw $21, 32($0)
    InstROM[13]  = 32'b00010010101101000000000000000011;             // beq $21, $20, 0x0003
    InstROM[14]  = 32'b10001100000101000000000000011111;             // lw $20, 31($0)
    InstROM[15]  = 32'b00010010101101000000000000000011;             // beq $21, $20, 0x0003
    InstROM[16]  = 32'b00000010010100011001100000100000;             // add $19, $18, $17
    InstROM[17]  = 32'b00000010001100001001000000100010;             // sub $18, $17, $16
    InstROM[18]  = 32'b00000010000011111000100000100011;             // subu $17, $16, $15
    InstROM[19]  = 32'b00001000000000000000000000001111;             // j 15
  end
  
endmodule

